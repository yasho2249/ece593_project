module rojo_module();


endmodule