// module rojo_tester(rojo_bfm bfm);


// endmodule: rojo_tester