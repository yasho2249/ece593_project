    Mac OS X            	   2  �     �                                    ATTR ��  �   �   �                  �   9  com.apple.quarantine        com.apple.lastuseddate#PS E5-  %   H  com.apple.macl 400081;61887da8;Chrome;E06E8400-3328-46E5-9C82-A5C837E2B441�߭a    �ud9     �2֟@��c���XT�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        This resource fork intentionally left blank                                                                                                                                                                                                                            ��